module dds(output reg [7:0] out,output reg sym,input [3:0] data,input wr,input clk);
reg [7:0] cos_list[0:255];
reg [7:0] cos_counter;
reg [3:0] split;
reg [3:0] split_count;
reg flag;

always @(negedge clk)
begin
	if(wr==1'b0)
	begin
	cos_counter<=8'h00;
	flag<=1'b0;
	sym<=1'b0;
	split<=data;
	split_count<=data;

	cos_list[0]<=8'hff;
	cos_list[1]<=8'hfe;
	cos_list[2]<=8'hfe;
	cos_list[3]<=8'hfe;
	cos_list[4]<=8'hfe;
	cos_list[5]<=8'hfe;
	cos_list[6]<=8'hfe;
	cos_list[7]<=8'hfe;
	cos_list[8]<=8'hfe;
	cos_list[9]<=8'hfe;
	cos_list[10]<=8'hfe;
	cos_list[11]<=8'hfe;
	cos_list[12]<=8'hfe;
	cos_list[13]<=8'hfe;
	cos_list[14]<=8'hfe;
	cos_list[15]<=8'hfd;
	cos_list[16]<=8'hfd;
	cos_list[17]<=8'hfd;
	cos_list[18]<=8'hfd;
	cos_list[19]<=8'hfd;
	cos_list[20]<=8'hfd;
	cos_list[21]<=8'hfc;
	cos_list[22]<=8'hfc;
	cos_list[23]<=8'hfc;
	cos_list[24]<=8'hfc;
	cos_list[25]<=8'hfb;
	cos_list[26]<=8'hfb;
	cos_list[27]<=8'hfb;
	cos_list[28]<=8'hfb;
	cos_list[29]<=8'hfa;
	cos_list[30]<=8'hfa;
	cos_list[31]<=8'hfa;
	cos_list[32]<=8'hfa;
	cos_list[33]<=8'hf9;
	cos_list[34]<=8'hf9;
	cos_list[35]<=8'hf9;
	cos_list[36]<=8'hf8;
	cos_list[37]<=8'hf8;
	cos_list[38]<=8'hf8;
	cos_list[39]<=8'hf7;
	cos_list[40]<=8'hf7;
	cos_list[41]<=8'hf6;
	cos_list[42]<=8'hf6;
	cos_list[43]<=8'hf6;
	cos_list[44]<=8'hf5;
	cos_list[45]<=8'hf5;
	cos_list[46]<=8'hf4;
	cos_list[47]<=8'hf4;
	cos_list[48]<=8'hf3;
	cos_list[49]<=8'hf3;
	cos_list[50]<=8'hf3;
	cos_list[51]<=8'hf2;
	cos_list[52]<=8'hf2;
	cos_list[53]<=8'hf1;
	cos_list[54]<=8'hf1;
	cos_list[55]<=8'hf0;
	cos_list[56]<=8'hef;
	cos_list[57]<=8'hef;
	cos_list[58]<=8'hee;
	cos_list[59]<=8'hee;
	cos_list[60]<=8'hed;
	cos_list[61]<=8'hed;
	cos_list[62]<=8'hec;
	cos_list[63]<=8'hec;
	cos_list[64]<=8'heb;
	cos_list[65]<=8'hea;
	cos_list[66]<=8'hea;
	cos_list[67]<=8'he9;
	cos_list[68]<=8'he8;
	cos_list[69]<=8'he8;
	cos_list[70]<=8'he7;
	cos_list[71]<=8'he6;
	cos_list[72]<=8'he6;
	cos_list[73]<=8'he5;
	cos_list[74]<=8'he4;
	cos_list[75]<=8'he4;
	cos_list[76]<=8'he3;
	cos_list[77]<=8'he2;
	cos_list[78]<=8'he2;
	cos_list[79]<=8'he1;
	cos_list[80]<=8'he0;
	cos_list[81]<=8'hdf;
	cos_list[82]<=8'hdf;
	cos_list[83]<=8'hde;
	cos_list[84]<=8'hdd;
	cos_list[85]<=8'hdc;
	cos_list[86]<=8'hdc;
	cos_list[87]<=8'hdb;
	cos_list[88]<=8'hda;
	cos_list[89]<=8'hd9;
	cos_list[90]<=8'hd8;
	cos_list[91]<=8'hd7;
	cos_list[92]<=8'hd7;
	cos_list[93]<=8'hd6;
	cos_list[94]<=8'hd5;
	cos_list[95]<=8'hd4;
	cos_list[96]<=8'hd3;
	cos_list[97]<=8'hd2;
	cos_list[98]<=8'hd1;
	cos_list[99]<=8'hd1;
	cos_list[100]<=8'hd0;
	cos_list[101]<=8'hcf;
	cos_list[102]<=8'hce;
	cos_list[103]<=8'hcd;
	cos_list[104]<=8'hcc;
	cos_list[105]<=8'hcb;
	cos_list[106]<=8'hca;
	cos_list[107]<=8'hc9;
	cos_list[108]<=8'hc8;
	cos_list[109]<=8'hc7;
	cos_list[110]<=8'hc6;
	cos_list[111]<=8'hc5;
	cos_list[112]<=8'hc4;
	cos_list[113]<=8'hc3;
	cos_list[114]<=8'hc2;
	cos_list[115]<=8'hc1;
	cos_list[116]<=8'hc0;
	cos_list[117]<=8'hbf;
	cos_list[118]<=8'hbe;
	cos_list[119]<=8'hbd;
	cos_list[120]<=8'hbc;
	cos_list[121]<=8'hbb;
	cos_list[122]<=8'hba;
	cos_list[123]<=8'hb9;
	cos_list[124]<=8'hb8;
	cos_list[125]<=8'hb7;
	cos_list[126]<=8'hb5;
	cos_list[127]<=8'hb4;
	cos_list[128]<=8'hb3;
	cos_list[129]<=8'hb2;
	cos_list[130]<=8'hb1;
	cos_list[131]<=8'hb0;
	cos_list[132]<=8'haf;
	cos_list[133]<=8'hae;
	cos_list[134]<=8'hac;
	cos_list[135]<=8'hab;
	cos_list[136]<=8'haa;
	cos_list[137]<=8'ha9;
	cos_list[138]<=8'ha8;
	cos_list[139]<=8'ha7;
	cos_list[140]<=8'ha5;
	cos_list[141]<=8'ha4;
	cos_list[142]<=8'ha3;
	cos_list[143]<=8'ha2;
	cos_list[144]<=8'ha1;
	cos_list[145]<=8'h9f;
	cos_list[146]<=8'h9e;
	cos_list[147]<=8'h9d;
	cos_list[148]<=8'h9c;
	cos_list[149]<=8'h9a;
	cos_list[150]<=8'h99;
	cos_list[151]<=8'h98;
	cos_list[152]<=8'h97;
	cos_list[153]<=8'h95;
	cos_list[154]<=8'h94;
	cos_list[155]<=8'h93;
	cos_list[156]<=8'h92;
	cos_list[157]<=8'h90;
	cos_list[158]<=8'h8f;
	cos_list[159]<=8'h8e;
	cos_list[160]<=8'h8c;
	cos_list[161]<=8'h8b;
	cos_list[162]<=8'h8a;
	cos_list[163]<=8'h88;
	cos_list[164]<=8'h87;
	cos_list[165]<=8'h86;
	cos_list[166]<=8'h84;
	cos_list[167]<=8'h83;
	cos_list[168]<=8'h82;
	cos_list[169]<=8'h80;
	cos_list[170]<=8'h7f;
	cos_list[171]<=8'h7e;
	cos_list[172]<=8'h7c;
	cos_list[173]<=8'h7b;
	cos_list[174]<=8'h7a;
	cos_list[175]<=8'h78;
	cos_list[176]<=8'h77;
	cos_list[177]<=8'h75;
	cos_list[178]<=8'h74;
	cos_list[179]<=8'h73;
	cos_list[180]<=8'h71;
	cos_list[181]<=8'h70;
	cos_list[182]<=8'h6e;
	cos_list[183]<=8'h6d;
	cos_list[184]<=8'h6c;
	cos_list[185]<=8'h6a;
	cos_list[186]<=8'h69;
	cos_list[187]<=8'h67;
	cos_list[188]<=8'h66;
	cos_list[189]<=8'h64;
	cos_list[190]<=8'h63;
	cos_list[191]<=8'h61;
	cos_list[192]<=8'h60;
	cos_list[193]<=8'h5f;
	cos_list[194]<=8'h5d;
	cos_list[195]<=8'h5c;
	cos_list[196]<=8'h5a;
	cos_list[197]<=8'h59;
	cos_list[198]<=8'h57;
	cos_list[199]<=8'h56;
	cos_list[200]<=8'h54;
	cos_list[201]<=8'h53;
	cos_list[202]<=8'h51;
	cos_list[203]<=8'h50;
	cos_list[204]<=8'h4e;
	cos_list[205]<=8'h4d;
	cos_list[206]<=8'h4b;
	cos_list[207]<=8'h4a;
	cos_list[208]<=8'h48;
	cos_list[209]<=8'h47;
	cos_list[210]<=8'h45;
	cos_list[211]<=8'h44;
	cos_list[212]<=8'h42;
	cos_list[213]<=8'h41;
	cos_list[214]<=8'h3f;
	cos_list[215]<=8'h3e;
	cos_list[216]<=8'h3c;
	cos_list[217]<=8'h3b;
	cos_list[218]<=8'h39;
	cos_list[219]<=8'h38;
	cos_list[220]<=8'h36;
	cos_list[221]<=8'h35;
	cos_list[222]<=8'h33;
	cos_list[223]<=8'h31;
	cos_list[224]<=8'h30;
	cos_list[225]<=8'h2e;
	cos_list[226]<=8'h2d;
	cos_list[227]<=8'h2b;
	cos_list[228]<=8'h2a;
	cos_list[229]<=8'h28;
	cos_list[230]<=8'h27;
	cos_list[231]<=8'h25;
	cos_list[232]<=8'h24;
	cos_list[233]<=8'h22;
	cos_list[234]<=8'h20;
	cos_list[235]<=8'h1f;
	cos_list[236]<=8'h1d;
	cos_list[237]<=8'h1c;
	cos_list[238]<=8'h1a;
	cos_list[239]<=8'h19;
	cos_list[240]<=8'h17;
	cos_list[241]<=8'h15;
	cos_list[242]<=8'h14;
	cos_list[243]<=8'h12;
	cos_list[244]<=8'h11;
	cos_list[245]<=8'hf;
	cos_list[246]<=8'he;
	cos_list[247]<=8'hc;
	cos_list[248]<=8'ha;
	cos_list[249]<=8'h9;
	cos_list[250]<=8'h7;
	cos_list[251]<=8'h6;
	cos_list[252]<=8'h4;
	cos_list[253]<=8'h3;
	cos_list[254]<=8'h1;
	cos_list[255]<=8'h0;
	end
	else
	begin
		if(split_count==split)
		begin
			out<=cos_list[cos_counter];
			if(flag==1'b0)cos_counter=cos_counter+1;
			else cos_counter=cos_counter-1;
			if(cos_counter==8'hfe)
			begin
				sym=~sym;
				flag=1'b1;
			end
			else if(cos_counter==8'h01)flag=1'b0;
			split_count<=4'b0000;
		end
		else
		begin
			split_count<=split_count+1;
		end
	end
end
endmodule
